`default_nettype none

module IzhilevichNeuron (


    
)